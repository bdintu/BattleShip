library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Joy is
	port(
		WASD : in std_logic_vector(4 downto 0)
	);
end Joy;

architecture Behavioral of Joy is
begin

end Behavioral;