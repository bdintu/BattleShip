library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity joy is
	port(
		WASD : in std_logic_vector(4 downto 0)
	);
end joy;

architecture Behavioral of joy is
begin

end Behavioral;